*
* ICL7652/101 OPERATIONAL AMPLIFIER "MACROMODEL" SUBCIRCUIT
* CREATED USING PARTS RELEASE 4.03 ON 08/07/90 AT 10:36
* REV (B)        SUPPLY VOLTAGE: +/-5V
* CONNECTIONS:   NON-INVERTING INPUT
*                | INVERTING INPUT
*                | | POSITIVE POWER SUPPLY
*                | | | NEGATIVE POWER SUPPLY
*                | | | | OUTPUT
*                | | | | |
.SUBCKT ICL7652/101_0   1 2 3 4 5
*
C1   11 12 3.804E-12
C2    6  7 20.00E-12
DC    5 53 DX
DE   54  5 DX
DLP  90 91 DX
DLN  92 90 DX
DP    4  3 DX
EGND 99  0 POLY(2) (3,0) (4,0) 0 .5 .5
FB 7 99 POLY(5) VB VC VE VLP VLN 0 1.342E9 -2E9 2E9 2E9 -2E9
GA    6  0 11 12 125.7E-6
GCM 0  6 10 99 25E-12
ISS   3 10 DC 56.00E-6
HLIM 90  0 VLIM 1K
J1   11  2 10 JX
J2   12  1 10 JX
R2    6  9 100.0E3
RD1 60 11 7.958E3
RD2 60 12 7.958E3
RO1   8  5 165
RO2   7 99 165
RP    3  4 6.667E3
RSS  10 99 3.571E6
VAD  60 4 -.7
VB    9  0 DC 0
VC 3 53 DC .84
VE   54  4 DC .74
VLIM  7  8 DC 0
VLP  91  0 DC 3.100
VLN   0 92 DC 3.100
.MODEL DX D(IS=800.0E-18)
.MODEL JX PJF(IS=500.0E-15 BETA=564.0E-6 VTO=-.183)
.ENDS
