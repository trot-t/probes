*
* OPA511 OPERATIONAL AMPLIFIER "MACROMODEL" SUBCIRCUIT
* "E" IS ENHANCED MODEL
* CREATED USING PARTS RELEASE 4.03 ON 09/11/90 AT 13:16
*
* REV.A 3/21/92 BCB: ADDED INPUT BIAS CURRENT CORRECTION
*
*
* CONNECTIONS:   NON-INVERTING INPUT
*                | INVERTING INPUT
*                | | POSITIVE POWER SUPPLY
*                | | | NEGATIVE POWER SUPPLY
*                | | | | OUTPUT
*                | | | | |
.SUBCKT OPA511_0   1 2 3 4 5
*
C1   11 12 20.00E-12
C2    6  7 40.00E-12
DC    5 53 DX
DE   54  5 DX
DLP  90 91 DX
DLN  92 90 DX
DP    4  3 DX
EGND 99  0 POLY(2) (3,0) (4,0) 0 .5 .5
FB    7 99 POLY(5) VB VC VE VLP VLN 0 8.950E9 -9E9 9E9 9E9 -9E9
GA    6  0 11 12 251.3E-6
GCM   0  6 10 99 794.8E-12
ISS   3 10 DC 160.0E-6
HLIM 90  0 VLIM 1K
J1   11  2 10 JX
J2   12  1 10 JX
G11 2 4 POLY(3) (10,2) (11,2) (4,2) 0 1E-12 1E-12 1E-12
G21 1 4 POLY(3) (10,1) (12,1) (4,1) 0 1E-12 1E-12 1E-12
R2    6  9 100.0E3
RD1   4 11 3.979E3
RD2   4 12 3.979E3
RO1   8  5 .25
RO2   7 99 .25
*  RP    3  4 2.800E3
RSS  10 99 1.250E6
VB    9  0 DC 0
VC    3 53 DC 5
VE   54  4 DC 5
VLIM  7  8 DC 0
VLP  91  0 DC 5.000E3
VLN   0 92 DC 5.000E3
****************************
* OPA511 "E" - ENHANCEMENTS
****************************
* OUTPUT SUPPLY MIRROR
FQ3   0 20 POLY(1) VLIM 0  1
DQ1  20 21 DX
DQ2  22 20 DX
VQ1  21  0 0
VQ2  22  0 0
FQ1   3  0 POLY(1) VQ1  19.62E-3  1
FQ2   0  4 POLY(1) VQ2  19.62E-3 -1
* QUIESCIENT CURRENT
RQ    3  4  2.5E5
* DIFF INPUT CAPACITANCE
CDIF  1  2  2.0E-12
* COMMON MODE INPUT CAPACITANCE
C1CM  1  99 2.0E-12
C2CM  2  99 2.0E-12
****************************
.MODEL DX D(IS=800.0E-18)
.MODEL JX PJF(IS=7.500E-9 BETA=197.4E-6 VTO=-1)
.ENDS
