*
* OP-07D/301 OPERATIONAL AMPLIFIER "MACROMODEL" SUBCIRCUIT
* CREATED USING PARTS RELEASE 4.01 ON 09/21/89 AT 09:26
* (REV N/A)      SUPPLY VOLTAGE: +/-15V
* CONNECTIONS:   NON-INVERTING INPUT
*                | INVERTING INPUT
*                | | POSITIVE POWER SUPPLY
*                | | | NEGATIVE POWER SUPPLY
*                | | | | OUTPUT
*                | | | | |
.SUBCKT OP-07D/301_0    1 2 3 4 5
*
C1   11 12 6.996E-12
C2    6  7 30.00E-12
DC    5 53 DX
DE   54  5 DX
DLP  90 91 DX
DLN  92 90 DX
DP    4  3 DX
EGND 99  0 POLY(2) (3,0) (4,0) 0 .5 .5
FB    7 99 POLY(5) VB VC VE VLP VLN 0 115.9E6 -100E6 100E6 100E6 -100E6
GA    6  0 11 12 115.0E-6
GCM   0  6 10 99 204.5E-12
IEE  10  4 DC 9.004E-6
HLIM 90  0 VLIM 1K
Q1   11  2 13 QX
Q2   12  1 14 QX
R2    6  9 100.0E3
RC1   3 11 8.696E3
RC2   3 12 8.696E3
RE1  13 10 2.947E3
RE2  14 10 2.947E3
REE  10 99 22.21E6
RO1   8  5 30
RO2 7 99 31.2
RP    3  4 11.29E3
VB    9  0 DC 0
VC    3 53 DC 2.800
VE   54  4 DC 2.800
VLIM  7  8 DC 0
VLP  91  0 DC 20
VLN   0 92 DC 20
.MODEL DX D(IS=800.0E-18)
.MODEL QX NPN(IS=800.0E-18 BF=2.250E3)
.ENDS
