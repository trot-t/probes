*//////////////////////////////////////////////////////////////////////
* (C) NATIONAL SEMICONDUCTOR, INC.
* MODELS DEVELOPED AND UNDER COPYRIGHT BY:
* NATIONAL SEMICONDUCTOR, INC.

*/////////////////////////////////////////////////////////////////////
* LEGAL NOTICE: THIS MATERIAL IS INTENDED FOR FREE SOFTWARE SUPPORT.
* THE FILE MAY BE COPIED, AND DISTRIBUTED; HOWEVER, RESELLING THE
*  MATERIAL IS ILLEGAL

*////////////////////////////////////////////////////////////////////
* FOR ORDERING OR TECHNICAL INFORMATION ON THESE MODELS, CONTACT:
* NATIONAL SEMICONDUCTOR'S CUSTOMER RESPONSE CENTER
*                 7:00 A.M.--7:00 P.M.  U.S. CENTRAL TIME
*                                (800) 272-9959
* FOR APPLICATIONS SUPPORT, CONTACT THE INTERNET ADDRESS:
*  AMPS-APPS@GALAXY.NSC.COM

*//////////////////////////////////////////////////////////
*LM741 OPERATIONAL AMPLIFIER MACRO-MODEL
*//////////////////////////////////////////////////////////
*
* CONNECTIONS:      NON-INVERTING INPUT
*                   |   INVERTING INPUT
*                   |   |   POSITIVE POWER SUPPLY
*                   |   |   |   NEGATIVE POWER SUPPLY
*                   |   |   |   |   OUTPUT
*                   |   |   |   |   |
*                   |   |   |   |   |
.SUBCKT LM741_0        1   2  99  50  28
*
* PINOUT ORDER +IN -IN V+ V- OUT
*
*
*FEATURES:
*IMPROVED PERFORMANCE OVER INDUSTRY STANDARDS
*PLUG-IN REPLACEMENT FOR LM709,LM201,MC1439,748
*INPUT AND OUTPUT OVERLOAD PROTECTION
*
****************INPUT STAGE**************
*
IOS 2 1 20N
*^INPUT OFFSET CURRENT
R1 1 3 250K
R2 3 2 250K
I1 4 50 100U
R3 5 99 517
R4 6 99 517
Q1 5 2 4 QX
Q2 6 7 4 QX
*FP2=2.55 MHZ
C4 5 6 60.3614P
*
***********COMMON MODE EFFECT***********
*
I2 99 50 1.6MA
*^QUIESCENT SUPPLY CURRENT
EOS 7 1 POLY(1) 16 49 1E-3 1
*INPUT OFFSET VOLTAGE.^
R8 99 49 40K
R9 49 50 40K
*
*********OUTPUT VOLTAGE LIMITING********
V2 99 8 1.63
D1 9 8 DX
D2 10 9 DX
V3 10 50 1.63
*
**************SECOND STAGE**************
*
EH 99 98 99 49 1
G1 98 9 5 6 2.1E-3
*FP1=5 HZ
R5 98 9 95.493MEG
C3 98 9 333.33P
*
***************POLE STAGE***************
*
*FP=30 MHZ
G3 98 15 9 49 1E-6
R12 98 15 1MEG
C5 98 15 5.3052E-15
*
*********COMMON-MODE ZERO STAGE*********
*
*FPCM=300 HZ
G4 98 16 3 49 3.1623E-8
L2 98 17 530.5M
R13 17 16 1K
*
**************OUTPUT STAGE**************
*
F6 50 99 POLY(1) V6 450U 1
E1 99 23 99 15 1
R16 24 23 25
D5 26 24 DX
V6 26 22 0.65V
R17 23 25 25
D6 25 27 DX
V7 22 27 0.65V
V5 22 21 0.18V
D4 21 15 DX
V4 20 22 0.18V
D3 15 20 DX
L3 22 28 100P
RL3 22 28 100K
*
***************MODELS USED**************
*
.MODEL DX D(IS=1E-15)
.MODEL QX NPN(BF=625)
*
.ENDS
