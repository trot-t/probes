* BEGIN MODEL LM7341
*//////////////////////////////////////////////////////////////////////
* (C) NATIONAL SEMICONDUCTOR, CORPORATION.
* MODELS DEVELOPED AND UNDER COPYRIGHT BY:
* NATIONAL SEMICONDUCTOR, CORPORATION.
*/////////////////////////////////////////////////////////////////////
* LEGAL NOTICE:
* THE MODEL MAY BE COPIED, AND DISTRIBUTED WITHOUT ANY MODIFICATIONS;
* HOWEVER, RESELLING OR LICENSING THE MATERIAL IS ILLEGAL.
* WE RESERVE THE RIGHT TO MAKE CHANGES TO THE MODEL WITHOUT PRIOR NOTICE.
* PSPICE MODELS ARE PROVIDED "AS IS, WITH NO WARRANTY OF ANY KIND"
*///////////////////////////////////////////////////////////////////
* PINOUT ORDER +IN -IN +V -V OUT
* PINOUT ORDER  3   4   5  2  1
.SUBCKT LM7341_0  3 4 5 2 1
*//////////////////////////////////////////
* SEE BELOW FOR PROGRAMMING INFORMATION
* SEE BELOW FOR MODEL FEATURES
* START PROGRAMMING
****************************
* BECAUSE THE PARAMETERS OF THE LM7341 VARY NOTICABLY AND NONLINEARLY
* WITH OPERATING VOLTAGE OVER THE WIDE OPERATING VOLTAGE RANGE OF THE
* PART (2.7 TO 30 VOLTS), THE MODEL IS PROGRAMMABLE TO SOME EXTENT.
* THERE ARE THREE GROUPS OF SPICE STATEMENTS FOR PROGRAMMING. ONLY
* ONE GROUP SHOULD BE UN-COMMENTED AT A TIME. THE THREE GROUPS ARE
* FOR 2.7, 10, AND 30 VOLTS TOTAL ACROSS THE PART. THE MODEL IS NOW
* SET UP FOR 10 VOLTS IE THE 10 VOLT GROUP IS UN-COMMENTED. FOR OTHER
* SUPPLY VOLTAGES THE VALUES MAY BE INTERPOLATED. SEE BELOW FOR AN
* INDEX TO THE FUNCTIONS OF THE PROGRAMMABLE COMPONENTS. V6 AND V7
* MAY BE ADJUSTED FOR ANY DESIRED OFFSET OR OFFSET DELTA FOR INPUT
* COMMON MODE NEAR THE POSITIVE RAIL.
************************************
* 2.7V GROUP
*V6 43 53 -350E-6
*V7 61 53 -10E-6
*G29 13 56 83 0 -7.5E-6
*R316 47 44 21
*R317 47 46 21
*R318 54 59 21
*R319 51 59 21
*R159 20 15 1.3E6
*E156 68 4 84 0 1.25
*E146 63 68 66 67 0.510
*G30 60 63 85 0 5E-6
*G27 60 63 64 65 8.5E-6
*I16 5 2 0.32E-3
*G25 5 2 42 0 0.3E-3
***************************************
* 10V GROUP
V6 43 53 -350E-6
V7 61 53 500E-6
G29 13 56 83 0 -8.5E-6
R316 47 44 19
R317 47 46 19
R318 54 59 19
R319 51 59 19
R159 20 15 2.7E6
E156 68 4 84 0 1.18
E146 63 68 66 67 0.335
G30 60 63 85 0 6.5E-6
G27 60 63 64 65 1E-5
I16 5 2 0.35E-3
G25 5 2 42 0 0.17E-3
******************************************
* 30V GROUP
*V6 43 53 -350E-6
*V7 61 53 1900E-6
*G29 13 56 83 0 -9.5E-6
*R316 47 44 15
*R317 47 46 15
*R318 54 59 15
*R319 51 59 15
*R159 20 15 6.0E6
*E156 68 4 84 0 1.04
*E146 63 68 66 67 0.345
*G30 60 63 85 0 6.5E-6
*G27 60 63 64 65 1E-5
*I16 5 2 0.41E-3
*G25 5 2 42 0 0.15E-3
**************************************
* END PROGRAMMING
* INDEX TO PROGRAMMABLE COMPONENT FUNCTIONS
* THE LINES IN THIS INDEX MUST ALWAYS REMAIN COMMENTED
*
*V6   RELATIVE OFFSET BETWEEN INPUT STAGES
*V7   OVERALL OFFSET
*G29  FRONT END CURRENT
*R316 BANDWIDTH/GAIN ADJ
*R317 BANDWIDTH/GAIN ADJ
*R318 BANDWIDTH/GAIN ADJ
*R319 BANDWIDTH/GAIN ADJ
*R159 DC GAIN ADJUST
*E156 VOLTAGE NOISE
*E146 VOLTAGE NOISE 1/F REGION
*G30  CURRENT NOISE
*G27  CURRENT NOISE 1/F REGION
*I16  IQ OFFSET
*G25  IQ TEMPERATURE SLOPE
*
* END OF INDEX
*///////////////////////////////////////////////
* MODEL FEATURES INCLUDE GAIN AND PHASE, SLEW RATE,
* VOLTAGE NOISE WITH 1/F, CURRENT NOISE WITH 1/F,
* INPUT BIAS CURRENT, INPUT BIAS CURRENT CHANGE
* WHEN COMMON MODE VOLTAGE NEAR THE + RAIL, INPUT
* OFFSET VOLTAGE, INPUT OFFSET VOLTAGE CHANGE WHEN
* WHEN COMMON MODE VOLTAGE NEAR THE + RAIL, INPUT
* OFFSET TEMPCO, COMMON MODE RANGE, CMRR WITH FREQ
* EFFECTS, PSRR WITH FREQ EFFECTS, OUTPUT SWING,
* OUTPUT CURRENT FLOWS THROUGH THE RAILS, OUTPUT
* CURRENT LIMIT, IQ AND IQ TEMPCO, AND CAPACATIVE
* LOAD EFFECTS.
*/////////////////////////////////////////////
Q41 6 7 8 QLN
R148 7 9 1E3
R149 10 11 1E3
R150 12 13 2.7
R151 8 14 2.7
R153 15 16 25
R154 17 13 2.7
R155 8 18 2.7
D22 19 5 DD
D23 2 19 DD
E58 8 0 2 0 1
E79 13 0 5 0 1
R156 2 5 1.1E9
E60 20 8 13 8 0.5
D24 21 13 DD
D25 8 22 DD
R157 23 24 100
R158 25 26 100
G14 15 20 27 20 0.1E-3
C24 16 28 15E-12
C25 19 0 0.5E-12
D26 26 6 DD
D27 29 24 DD
Q42 29 11 13 QLP
R160 19 30 1
R161 31 19 1
E71 32 20 33 34 -1
R162 32 27 1E4
C26 27 20 0.3E-12
G15 35 20 15 20 -1E-3
G16 20 36 15 20 1E-3
G17 20 37 38 8 1E-3
G18 39 20 13 40 1E-3
D28 39 35 DD
D29 36 37 DD
R163 35 39 1E9
R164 37 36 1E9
R165 39 13 1E3
R166 8 37 1E3
R167 36 20 1E7
R168 37 20 1E7
R169 20 39 1E7
R170 20 35 1E7
R171 20 27 1E9
R172 23 13 1E9
R173 8 25 1E9
G20 40 38 41 0 0.3E-3
L2 19 1 0.4E-9
R175 19 1 4E2
R176 40 13 1E8
R177 8 38 1E8
R178 14 26 1E8
R179 12 24 1E8
E84 13 10 13 12 9
E85 9 8 14 8 9
E24 28 0 19 0 1
R219 15 28 6E8
Q52 30 24 12 QOP
Q53 31 26 14 QON
Q54 38 38 18 QON
Q55 40 40 17 QOP
E144 13 23 13 39 1
E145 25 8 37 8 1
E51 15 22 20 8 0.7
E52 21 15 13 20 0.7
G23 5 0 30 19 1
G24 2 0 19 31 -1
Q56 33 43 44 QIN
Q57 34 45 46 QIN
Q58 47 48 8 Q
Q59 48 49 8 Q
Q60 50 45 51 QIP
Q61 52 53 54 QIP
Q62 55 56 13 QP
Q63 48 57 58 QPX
R320 60 61 200
R321 33 13 300
R322 8 50 300
R323 8 52 300
V4 13 62 1
R324 63 45 200
D30 43 13 DD
D31 45 13 DD
D32 8 53 DD
D33 8 45 DD
D34 64 0 DIN
D35 65 0 DIN
I9 0 64 0.1E-3
I10 0 65 0.1E-3
C27 60 0 1E-12
C28 4 0 1E-12
D36 66 0 DVN
D37 67 0 DVN
I11 0 66 0.1E-3
I12 0 67 0.1E-3
E147 69 0 13 0 1
E148 70 0 8 0 1
E149 71 0 72 0 1
R329 69 73 1E6
R330 70 74 1E6
R331 71 75 1E6
R332 0 73 100
R333 0 74 100
R334 0 75 1E4
E150 76 3 75 0 1E-6
R335 63 72 1E9
R336 72 60 1E9
C29 69 73 1E-12
C30 70 74 3E-12
C31 71 75 1E-12
R337 34 13 300
E151 77 76 74 0 -0.7
E152 78 77 73 0 0.7
C32 34 33 4E-12
C33 50 52 4E-12
G28 15 20 79 20 0.1E-3
E153 80 20 50 52 1
R338 80 79 1E4
C34 79 20 0.3E-12
R339 20 79 1E9
V12 41 0 1
V15 55 59 0
R341 55 58 1
R342 57 62 1E4
R343 48 49 80
I14 0 81 1E-3
D39 81 0 DD
R345 0 82 1E7
E155 83 0 82 0 -1.75
R346 0 83 1E7
V17 81 82 1.2301
R347 0 84 9.6E4
R348 0 84 9.6E4
R349 0 85 9.6E4
R350 0 85 9.6E4
E158 60 78 42 0 1.125E-3
I15 0 86 1E-3
D40 86 0 DD
R352 0 42 1E7
V19 86 42 0.655
R353 78 60 1E9
R354 77 78 1E9
R355 76 77 1E9
R356 3 76 1E9
R357 0 41 1E9
.MODEL QON NPN RC=1 IS=1E-13
.MODEL QOP PNP RC=1 IS=1E-13
.MODEL QPX PNP BF=200 IS=1E-14
.MODEL DD D
.MODEL QIN NPN BF=1.2E4
.MODEL QIP PNP BF=4.4E3
.MODEL Q NPN
.MODEL QP PNP
.MODEL DVN D KF=2.5E-15
.MODEL DIN D KF=1E-15
.MODEL QLN NPN
.MODEL QLP PNP
.ENDS
