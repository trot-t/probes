title
* комментарий
XU1 1 3 plus minus 5 LF356_0
R3 1 0 1k
R1 2 1 1k
R2 3 4 1k
R4 3 5 1k
V1 2 0 0.1v  ; входной сигнал
V2 4 0 0v  

.include 'LF356.cir'  ; подключить файл со схемой операционного усилителя

Vplus plus 0 15     ; питание микросхемы
Vminus 0 minus 15   ; питание микросхемы

.control
set color0 = white  ; пожалеть принтер, цвет фона - белый
*tran 0.1m 1        ; анализ переходных процессов
DC V1 0 20 0.1      ; анализ при постоянном токе
plot v(5)    ; график выходного сигнала
* если есть gnuplot график будет выведен в файл how_to_use.png (если нет gnuplot, файл с графиком не создастся, ошибки не повлияют на выполнение)
set gnuplot_terminal=png/quit
gnuplot  how_to_use v(5)
.endc

.end
