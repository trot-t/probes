* OPA445E OPERATIONAL AMPLIFIER "MACROMODEL" SUBCIRCUIT
* CREATED USING PARTS RELEASE 4.03 ON 10/04/90 AT 14:31
*
* REV.B 3/21/92 BCB: ADDING INPUT BIAS CURRENT CORRECTION
*
* ------------------------------------------------------------------------
*|(C) COPYRIGHT TEXAS INSTRUMENTS INCORPORATED 2007. ALL RIGHTS RESERVED. |
*|                                                                        |
*|THIS MODEL IS DESIGNED AS AN AID FOR CUSTOMERS OF TEXAS INSTRUMENTS.    |
*|NO WARRANTIES, EITHER EXPRESSED OR IMPLIED, WITH RESPECT TO THIS MODEL  |
*|OR ITS FITNESS FOR A PARTICULAR PURPOSE IS CLAIMED BY TEXAS INSTRUMENTS |
*|OR THE AUTHOR.  THE MODEL IS LICENSED SOLELY ON AN "AS IS" BASIS.  THE  |
*|ENTIRE RISK AS TO ITS QUALITY AND PERFORMANCE IS WITH THE CUSTOMER.     |
* ------------------------------------------------------------------------
*
* CONNECTIONS:   NON-INVERTING INPUT
*                | INVERTING INPUT
*                | | POSITIVE POWER SUPPLY
*                | | | NEGATIVE POWER SUPPLY
*                | | | | OUTPUT
*                | | | | |
.SUBCKT OPA445E_0   1 2 3 4 5
*
C1   11 12 5.252E-12
C2    6  7 15.00E-12
DC    5 53 DX
DE   54  5 DX
DLP  90 91 DX
DLN  92 90 DX
DP    4  3 DX
EGND 99  0 POLY(2) (3,0) (4,0) 0 .5 .5
FB    7 99 POLY(5) VB VC VE VLP VLN 0 37.74E6 -40E6 40E6 40E6 -40E6
GA    6  0 11 12 188.5E-6
GCM   0  6 10 99 3.352E-9
ISS   3 10 DC 202.5E-6
HLIM 90  0 VLIM 1K
J1   11  2 10 JX
J2   12  1 10 JX
G11 2 4 POLY(3) (10,2) (11,2) (4,2) 0 1E-12 1E-12 1E-12
G21 1 4 POLY(3) (10,1) (12,1) (4,1) 0 1E-12 1E-12 1E-12
R2    6  9 100.0E3
RD1   4 11 5.305E3
RD2   4 12 5.305E3
RO1   8  5 25
RO2   7 99 25
*  RP    3  4 21.05E3
RSS  10 99 987.7E3
VB    9  0 DC 0
VC    3 53 DC 5
VE   54  4 DC 5
VLIM  7  8 DC 0
VLP  91  0 DC 26
VLN   0 92 DC 26
****************************
* OPA445 "E" - ENHANCEMENTS
****************************
* OUTPUT SUPPLY MIRROR
FQ3   0 20 POLY(1) VLIM 0  1
DQ1  20 21 DX
DQ2  22 20 DX
VQ1  21  0 0
VQ2  22  0 0
FQ1   3  0 POLY(1) VQ1  2.795E-3  1
FQ2   0  4 POLY(1) VQ2  2.795E-3 -1
* QUIESCIENT CURRENT
RQ    3  4  1.0E5
* DIFF INPUT CAPACITANCE
CDIF  1  2  1.0E-12
* COMMON MODE INPUT CAPACITANCE
C1CM  1  99 1.5E-12
C2CM  2  99 1.5E-12
****************************
.MODEL DX D(IS=800.0E-18)
.MODEL JX PJF(IS=10.00E-12 BETA=87.73E-6 VTO=-1)
.ENDS
