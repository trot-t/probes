*
* LT1013/5_1 OPERATIONAL AMPLIFIER "MACROMODEL" SUBCIRCUIT
* CREATED USING PARTS RELEASE 4.03 ON 07/18/90 AT 11:04
* REV (N/A)      SUPPLY VOLTAGE: 5V
* CONNECTIONS:   NON-INVERTING INPUT
*                | INVERTING INPUT
*                | | POSITIVE POWER SUPPLY
*                | | | NEGATIVE POWER SUPPLY
*                | | | | OUTPUT
*                | | | | |
.SUBCKT LT1013/5_1_0    1 2 3 4 5
*
C1   11 12 5.887E-12
C2    6  7 30.00E-12
DC    5 53 DX
DE   54  5 DX
DLP  90 91 DX
DLN  92 90 DX
DP    4  3 DX
EGND 99  0 POLY(2) (3,0) (4,0) 0 .5 .5
FB 7 99 POLY(5) VB VC VE VLP VLN 0 204.6E6 -20E6 20E6 20E6 -20E6
GA    6  0 11 12 113.1E-6
GCM   0  6 10 99 225.7E-12
IEE   3 10 DC 12.04E-6
HLIM 90  0 VLIM 1K
Q1   11  2 13 QX
Q2   12  1 14 QX
R2    6  9 100.0E3
RC1   4 11 8.842E3
RC2   4 12 8.842E3
RE1  13 10 4.518E3
RE2  14 10 4.518E3
REE  10 99 16.62E6
RO1   8  5 25
RO2   7 99 50
RP    3  4 16.23E3
VB    9  0 DC 0
VC    3 53 DC 1.300
VE   54  4 DC .7
VLIM  7  8 DC 0
VLP  91  0 DC 25
VLN   0 92 DC 25
.MODEL DX D(IS=800.0E-18)
.MODEL QX PNP(IS=800.0E-18 BF=333.3)
.ENDS
