* TLC2654 OPERATIONAL AMPLIFIER "MACROMODEL" SUBCIRCUIT
* CREATED USING PARTS RELEASE 4.03 ON 06/26/90 AT 08:49
* REV (N/A)      SUPPLY VOLTAGE: +/-5V  
* ------------------------------------------------------------------------
*|(C) COPYRIGHT TEXAS INSTRUMENTS INCORPORATED 2007. ALL RIGHTS RESERVED. |
*|                                                                        |
*|THIS MODEL IS DESIGNED AS AN AID FOR CUSTOMERS OF TEXAS INSTRUMENTS.    |
*|NO WARRANTIES, EITHER EXPRESSED OR IMPLIED, WITH RESPECT TO THIS MODEL  |
*|OR ITS FITNESS FOR A PARTICULAR PURPOSE IS CLAIMED BY TEXAS INSTRUMENTS |
*|OR THE AUTHOR.  THE MODEL IS LICENSED SOLELY ON AN "AS IS" BASIS.  THE  |
*|ENTIRE RISK AS TO ITS QUALITY AND PERFORMANCE IS WITH THE CUSTOMER.     |
* ------------------------------------------------------------------------
* CONNECTIONS:   NON-INVERTING INPUT
*                | INVERTING INPUT
*                | | POSITIVE POWER SUPPLY
*                | | | NEGATIVE POWER SUPPLY
*                | | | | OUTPUT
*                | | | | |
.SUBCKT TLC2654_0   1 2 3 4 5
*
C1   11 12 4.004E-12
C2    6  7 20.00E-12
C3   87 0 19.8E-9
CPSR 85 86 15.9E-6
DCM+ 81 82 DX
DCM- 83 81 DX
DC    5 53 DX
DE   54  5 DX
DLP  90 91 DX
DLN  92 90 DX
DP    4  3 DX
ECMR 84 99 (2,99) 1
EGND 99  0 POLY(2) (3,0) (4,0) 0 .5 .5
EPSR 85 0 POLY(1) (3,4) -22.7E-6  2.27E-6
ENSE 89 2 POLY(1) (88,0) 5E-6 1
FB 7 99 POLY(6) VB VC VE VLP VLN VPSR 0 1.798E9 -1E9 1E9 1E9 -1E9 1.236E9
GA    6  0 11 12 138.2E-6
GCM 0  6 10 99 154.73E-12
GPSR 85 86 (85,86) 100E-6
GRD1 60 11 (60,11) 1.382E-4
GRD2 60 12 (60,12) 1.382E-4
HLIM 90  0 VLIM 1K
HCMR 80 1 POLY(2) VCM+ VCM- 0 1E2 1E2
IRP 3 4 1.46E-3
ISS   3 10 DC 40.00E-6
IIO 2 0 30E-12
I1 88 0 1E-21
J1   11  89 10 JX
J2   12  80 10 JX
R2    6  9 100.0E3
RCM 84 81 1K
RN1 87 0 134E3
RN2 87 88 5E3
RO1   8  5 165
RO2   7 99 165
RSS  10 99 5.000E6
VAD  60 4 -.4
VCM+ 82 99 2.3
VCM- 83 99 -4.6
VB    9  0 DC 0
VC    3 53 DC .9
VE   54  4 DC .8
VLIM  7  8 DC 0
VLP  91  0 DC 3.100
VLN   0 92 DC 3.100
VPSR 0 86 DC 0
.MODEL DX D(IS=800.0E-18)
.MODEL JX PJF(IS=25.00E
