*//////////////////////////////////////////////////////////////////////
* (C) NATIONAL SEMICONDUCTOR, INC.
* MODELS DEVELOPED AND UNDER COPYRIGHT BY:
* NATIONAL SEMICONDUCTOR, INC.

*/////////////////////////////////////////////////////////////////////
* LEGAL NOTICE: THIS MATERIAL IS INTENDED FOR FREE SOFTWARE SUPPORT.
* THE FILE MAY BE COPIED, AND DISTRIBUTED; HOWEVER, RESELLING THE
*  MATERIAL IS ILLEGAL

*////////////////////////////////////////////////////////////////////
* FOR ORDERING OR TECHNICAL INFORMATION ON THESE MODELS, CONTACT:
* NATIONAL SEMICONDUCTOR'S CUSTOMER RESPONSE CENTER
*                 7:00 A.M.--7:00 P.M.  U.S. CENTRAL TIME
*                                (800) 272-9959
* FOR APPLICATIONS SUPPORT, CONTACT THE INTERNET ADDRESS:
*  AMPS-APPS@GALAXY.NSC.COM

* //////////////////////////////////////////
* LM4250 PROGRAMMABLE OPERATIONAL AMPLIFIER
* //////////////////////////////////////////
*
* CONNECTIONS:      NON-INVERTING INPUT
*                   |   INVERTING INPUT
*                   |   |   POSITIVE POWER SUPPLY
*                   |   |   |   NEGATIVE POWER SUPPLY
*                   |   |   |   |   OUTPUT
*                   |   |   |   |   |   QUIESCENT CURRENT SET
*                   |   |   |   |   |   |
.SUBCKT LM4250_0       3   2   6   4   7   8
*
* PINOUT ORDER +IN -IN V+ V- OUT SET
*
*
* FEATURES:
* +/-1V TO +/-18V POWER SUPPLY OPERATION
* INPUT OFFSET CURRENT (ISET=1UA) =      3NA
* LOW OFFSET VOLTAGE (TYP) =             2MV
* SLEW RATE =                         .2V/US
* GAIN-BANDWIDTH PRODUCT =            230KHZ
* MAX SUPPLY CURRENT (ISET=10UA) =     100UA
* SHORT CIRCUIT PROTECTED
*
* NOTE: - NOISE IS NOT MODELED.
*       - ASYMMETRICAL GAIN IS NOT MODELED.
*
* INPUT CAPACITORS.
CI1   3  4  2P
CI2   2  4  2P
* PRIMARY POLE=939.2MHZ.
C3    98 20 169.3N
* SECONDARY POLE=276KHZ.
C4    13 14 75.3P
C6    4  9  3P
* THIRD POLE=795KHZ.
C7    98 19 200E-15
D1    10 8  DX
D2    7  6  DX
D3    4  7  DX
D4    4  26 DX
D5    26 7  DX
D6    20 24 DX
D7    25 20 DX
D8    22 0  DX
D9    0  21 DX
D10   7  27 DX
D11   27 6  DX
* DETERMINES DC CMRR.
ECMRR 1  3  16        49 1.0
EH    97 98 6         49 1.0
EN    0  96 0         4  1.0
EP    97 0  6         0  1.0
E1    97 18 6         19 1.0
F1    6  0  VA2       1
F2    0  4  VA3       1
F3    23 0  VA1       1
F4    6  9  V1        1.0
F5    6  4  POLY(2)   V1 V5 0 8.0 0 0 1
* SETS -ISC
F6    4 26  POLY(1)   VA1 -1E-2 -1
* SETS +ISC
F7    27 6  POLY(1)   VA1 -1.2E-2 1
G1    98 20 14        13 1.0
G2    98 19 20        49 1U
G4    98 16 POLY(2) 3 49 2 49 0 1.581E-7 1.581E-7
G5    15 4  6         4  0.0333
* CMRR ZERO.
L2    16 17 73.1M
* IS OF QX1/QX2 AND R1/R2 DETERMINES VOS.
Q1    13 1  11        QX1
Q2    14 2  12        QX2
R1    9  11 9.6K
R2    9  12 10K
R3    14 4  3.83K
R4    13 4  3.83K
R5    98 20 1E6
R8    6  49 1E8
R9    49 4  1E8
R12   98 19 1E6
R13   98 17 1K
* OUTPUT RESISTANCE.
R22   28 7  581
VA1   18 28 0V
VA2   21 23 0V
VA3   23 22 0V
V1    6  10 0V
V2    97 24 1.5V
V3    25 96 1.5V
V5    4  15 0V
.MODEL QX1 PNP (IS=4.625E-16 BF=270 VAF=60 IKF=1E-3 NE=1.15 ISE=.63E-16)
.MODEL QX2 PNP (IS=5E-16 BF=300 VAF=60 IKF=1E-3 NE=1.15 ISE=.63E-16)
.MODEL DX D(IS=5E-15)
.ENDS
